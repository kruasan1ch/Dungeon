0;Am Shegar;1;117;erdwsgf
2;aesdfaw;1;130;vxc b
1;sfasdg;1;130;azdvs
0;Am Shegar;1;117;wadsd
2;aeega;1;130;awdsawfa
0;Am Shegar;1;117;awdasd
0;Am Shegar;1;117;awsdawd
0;awdfadf;1;117;awdas
0;123;1;117;124w4
0;Am Shegar;1;117;adsf
0;Am Shegar;1;117;sfgevsag
0;AWFAwf;1;117;adsawd

0;62;62;3;10;1;10;Am Shegar;1;117;150;5
0;45;65;3;20;1;20;Am Shegar;3;157;225;8